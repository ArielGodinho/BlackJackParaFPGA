library ieee;
use ieee.std_logic_1164.all;

entity Deck is
	port(
	);
end Deck;

architecture arch of Deck is
begin

end arch;