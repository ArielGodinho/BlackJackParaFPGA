library ieee;
use ieee.std_logic_1164.all;

entity Blackjack is
	port(
	);
end Blackjack;

architecture arch of Blackjack is

	signal 

begin

end arch;