library ieee;
use ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity TopLevelEntity is
	port(
		clock                : in  std_logic;
		reset                : in  std_logic
	);
end TopLevelEntity;

architecture arch of TopLevelEntity is
	
begin

end arch;
