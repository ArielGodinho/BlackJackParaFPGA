library ieee;
use ieee.std_logic_1164.all;

entity ControlUnit is
	port(
	);
end ControlUnit;

architecture arch of ControlUnit is

	signal 

begin
	process ()
	begin

	end process;

end arch ; -- archControlUnit