library ieee;
use ieee.std_logic_1164.all;

entity ResultCalculator is
	port(
	);
end ResultCalculator;

architecture arch of ResultCalculator is

	signal 

begin

end arch;