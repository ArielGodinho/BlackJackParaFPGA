library ieee;
use ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity TerminalInterface is
	port(
		clock                : in  std_logic;
		reset                : in  std_logic
	);
end TerminalInterface;

architecture arch of TerminalInterface is
	
begin

end arch;
